*   BF862 SPICE MODEL MARCH 2007 NXP SEMICONDUCTORS
*   ENVELOPE    SOT23
*   JBF862: 1, Drain,  2,Gate,  3,Source
.SUBCKT BF862 1 2 3
  Ld  1 4  L=	1.1nH
  Ls  3 6  L=	1.25nH
  Lg  2 5  L=	0.78nH
  Rg  5 7  R=	0.535 Ohm
  Cds  1 3  C=	0.0001pF
  Cgs  2 3  C=	1.05pF
  Cgd  1 2  C=	0.201pF
  Co  4 6  C=	0.35092pF
  Q1 4 7 6 JBF862
.model JBF862 NJF(Beta=47.800E-3 Betatce=-.5 Rd=.8 Rs=7.5000 Lambda=37.300E-3 Vto=-.57093
+ Vtotc=-2.0000E-3 Is=424.60E-12 Isr=2.995p N=1 Nr=2 Xti=3 Alpha=-1.0000E-3
+ Vk=59.97 Cgd=7.4002E-12 M=.6015 Pb=.5 Fc=.5 Cgs=8.2890E-12 Kf=87.5E-18
+ Af=1)
.ENDS BF862